module Bus#(
	int NUMBER_OF_CACHES = 4
)();
endmodule : Bus
