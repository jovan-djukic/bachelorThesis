package MSIStates;
	typedef enum logic[1 : 0] {
		INVALID,
		SHARED,
	  MODIFIED	
	} CacheLineState;
endpackage : MSIStates
