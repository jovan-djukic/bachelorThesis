package states;
	typedef enum logic[1 : 0] {
		INVALID,
		VALID,
		DIRTY
	} CacheLineState;
endpackage : states
